module top_module( output one );

// Insert your code hereassign one = 1'b1;
	
endmodule
