module top_module( 
  input x3,
  input x2,
  input x1,  // three inputs
  output f   // one output
);

endmodule